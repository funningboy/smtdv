
// 4x4 bus Matrix
