
`ifndef __APB_SLAVE_VSEQS_LIB_SV__
`define __APB_SLAVE_VSEQS_LIB_SV__

`include "apb_slave_base_vseq.sv"

`endif //__APB_SLAVE_VSEQS_LIB_SV__

