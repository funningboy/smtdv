
`ifndef __SMTDV_MODEL_LIB_SV__
`define __SMTDV_MODEL_LIB_SV__

`include "smtdv_generic_memory_cb.sv"
`include "smtdv_generic_memory.sv"
`include "smtdv_generic_fifo_cb.sv"
`include "smtdv_generic_fifo.sv"
`include "smtdv_ring_queue.sv"
`include "smtdv_reset_model.sv"
`include "smtdv_reset_monitor.sv"

// `include "smtdv_arbiter.sv"
// `include "smtdv_multi2one_channels.sv"
// `include "smtdv_one2multi_channels.sv"
// `include "smtdv_lowpower_model.sv"
// `include "ssmtdv_jtag_model.sv"

`endif // __SMTDV_MODEL_LIB_SV__
