
`ifndef __APB_FWCTRL_TEST_SV__
`define __APB_FWCTRL_TEST_SV__





`endif // end of __APB_FWCTRL_TEST_SV__
