../../../../../../../adapters/uvm_sv/uvm_ml_adapter_imp.sv