../../../../../../../adapters/uvm_sv/uvm_ml_phase_participate_handler.svh