`ifndef __AHB_TEST_LIST_SV__
`define __AHB_TEST_LIST_SV__

`timescale 1ns/10ps

package test_ahb_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import smtdv_sqlite3_pkg::*;
  import smtdv_stl_pkg::*;

  import smtdv_common_pkg::*;
  `include "smtdv_macros.svh"

  `include "ahb_defines.svh"
  import ahb_pkg::*;
  import ahb_seq_pkg::*;

`include "ahb_base_test.sv"
`include "ahb_setup_test.sv"
`include "ahb_rand_test.sv"
`include "ahb_stl_test.sv"
`include "ahb_busy_test.sv"
`include "ahb_split_test.sv"
`include "ahb_retry_test.sv"
`include "ahb_err_inject_test.sv"
`include "ahb_hijack_test.sv"
`include "ahb_polling_test.sv"
`include "ahb_interrupt_test.sv"
`include "ahb_incr_test.sv"
`include "ahb_swap_test.sv"
`include "ahb_wrap_test.sv"
//`include "ahb_fw_ctl_test.sv"
//`include "ahb_csim_test.sv"

endpackage

`endif // end of __AHB_TEST_LIST_SV__
