    class bogus;
    endclass
