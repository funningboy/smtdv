
`ifndef __SMTDV_LIB_SV__
`define __SMTDV_LIB_SV__

`include "smtdv_lib_typedefs.svh"
`include "smtdv_lib_utils.sv"
`include "smtdv_queue.sv"
`include "smtdv_hash.sv"
`include "smtdv_sequence.sv"
`include "smtdv_sequence_item.sv"
`include "smtdv_sequence_frame.sv"
`include "smtdv_component.sv"
`include "smtdv_cfg.sv"
`include "smtdv_slave_cfg.sv"
`include "smtdv_master_cfg.sv"
`include "smtdv_label.sv"
`include "smtdv_cfg_label.sv"
`include "smtdv_force_vif_label.sv"
`include "smtdv_force_block_label.sv"
`include "smtdv_force_rsp_err_label.sv"
`include "smtdv_force_replay_label.sv"
`include "smtdv_system_table.sv"
`include "smtdv_label_handler.sv"
`include "smtdv_thread.sv"
`include "smtdv_thread_handler.sv"
`include "smtdv_sequencer.sv"
`include "smtdv_push_sequencer.sv"
`include "smtdv_force_vif_threads.sv"
`include "smtdv_rsp_back_threads.sv"
`include "smtdv_ready_notify_threads.sv"
//`include "smtdv_lock_notify_threads.sv"
`include "smtdv_driver.sv"
`include "smtdv_push_driver.sv"
`include "smtdv_monitor.sv"
`include "smtdv_agent.sv"
`include "smtdv_master_agent.sv"
`include "smtdv_slave_agent.sv"
`include "smtdv_backdoor_threads.sv"
`include "smtdv_mem_bkdor_wr_cmp_threads.sv"
`include "smtdv_mem_bkdor_rd_cmp_threads.sv"
`include "smtdv_backdoor.sv"
`include "smtdv_scoreboard_threads.sv"
`include "smtdv_scoreboard_wr_threads.sv"
`include "smtdv_scoreboard_rd_threads.sv"
`include "smtdv_scoreboard.sv"
`include "smtdv_test.sv"
`include "smtdv_runtime_phases.svh"
`include "smtdv_report_server.sv"
`include "smtdv_reg_adapter.sv"

`endif
