// detect deadlock threads and kill
//
