`ifndef __UART_TYPEDEFS_SV__
`define __UART_TYPEDEFS_SV__

typedef enum bit {GOOD_PARITY, BAD_PARITY} parity_e;

`endif // __UART_TYPEDEFS_SV__
