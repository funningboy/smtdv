
`ifndef __APB_TEST_PKG_SV__
`define __APB_TEST_PKG_SV__

`timescale 1ns/10ps

package test_apb_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import smtdv_sqlite3_pkg::*;
  import smtdv_stl_pkg::*;

  import smtdv_common_pkg::*;
  `include "smtdv_macros.svh"

  `include "apb_defines.svh"
  `include "apb_macros.svh"

  import apb_pkg::*;
  import apb_seq_pkg::*;
  import apb_vseq_pkg::*;

  `include "apb_test_lib.sv"

endpackage : test_apb_pkg

`endif // end of __APB_TEST_PKG_SV__
