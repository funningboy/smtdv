`ifndef __AHB_PKG_SV__
`define __AHB_PKG_SV__

package ahb_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import smtdv_common_pkg::*;
  `include "smtdv_macros.svh"

  import smtdv_sqlite3_pkg::*;

  import smtdv_stl_pkg::*;

  `include "ahb_typedefs.svh"
  `include "ahb_item.sv"

  `include "ahb_monitor_threads.sv"
  `include "ahb_monitor.sv"

  `include "ahb_master_cfg.sv"
  `include "ahb_master_driver_threads.sv"
  `include "ahb_master_driver.sv"
  `include "ahb_master_sequencer.sv"
  `include "ahb_master_agent.sv"

  `include "ahb_slave_cfg.sv"
  `include "ahb_slave_driver_threads.sv"
  `include "ahb_slave_driver.sv"
  `include "ahb_slave_sequencer.sv"
  `include "ahb_slave_agent.sv"

  `include "ahb_scoreboard.sv"
  `include "ahb_reg_adapter.sv"

endpackage : ahb_pkg

`include "ahb_if.sv"

`endif
