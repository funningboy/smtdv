`ifndef __APB_TEST_LIST_SV__
`define __APB_TEST_LIST_SV__

`include "apb_base_env.sv"
`include "apb_base_test.sv"

`include "apb_setup_test.sv"
`include "apb_stl_test.sv"
`include "apb_err_inject_test.sv"
`include "apb_hijack_test.sv"
`include "apb_polling_test.sv"
`include "apb_interrupt_test.sv"
`include "apb_cfg_label_test.sv"
`include "apb_rand_test.sv"
`include "apb_csim_test.sv"

`endif // __APB_TEST_LIST_SV__
