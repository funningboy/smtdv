`ifndef __APB_TYPEDEFS_SV__
`define __APB_TYPEDEFS_SV__

typedef enum bit [0:0] {OK, ERR} trx_rsp_t;

`endif
