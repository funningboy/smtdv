
`ifndef __APB_SLAVE_SEQS_LIB_SV__
`define __APB_SLAVE_SEQS_LIB_SV__

`include "apb_slave_base_seq.sv"
`include "apb_slave_seqs.sv"
`include "apb_slave_err_inject_seq.sv"
`include "apb_slave_hijack_seq.sv"

`endif // __APB_SLAVE_SEQS_LIB_SV__
