
`ifndef __SMTDV_MASTER_SEQS_LIB_SV__
`define __SMTDV_MASTER_SEQS_LIB_SV__

`include "smtdv_master_base_seq.sv"
`include "smtdv_master_retry_seq.sv"
`include "smtdv_master_polling_seq.sv"
`include "smtdv_master_stop_seqr_seq.sv"
`include "smtdv_master_dump_memreg_seq.sv"
`include "smtdv_master_test_seq.sv"

`endif // __SMTDseqrseqr_
