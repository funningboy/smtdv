`ifndef __AHB_MASTER_VSEQS_LIB_SV__
`define __AHB_MASTER_VSEQS_LIB_SV__

`include "ahb_master_base_vseq.sv"
`include "ahb_master_1w1r_vseq.sv"
`include "ahb_master_rand_vseq.sv"
`include "ahb_master_retry_vseq.sv"
`include "ahb_master_polling_vseq.sv"
`include "ahb_master_interrupt_vseq.sv"
`include "ahb_master_mutex_vseq.sv"
`include "ahb_master_fw_ctl_vseq.sv"
//`include "ahb_master_reg_cfg_vseq.sv"

`endif // __AHB_MASTER_VSEQS_LIB_SV__
