
/*
*  declare all type of seqs
*/

`ifdef SMTDV_SEQ_32X32
    `SMTDV_MAGIC_SEQ_DEC(smtdv, 32, 32)
`endif

`ifdef SMTDV_SEQ_64X64
    `SMTDV_MAGIC_SEQ_DEC(smtdv, 64, 64)
`endif

