
`ifndef __SMTDV_LIB_SV__
`define __SMTDV_LIB_SV__

`include "smtdv_lib_typedefs.svh"
`include "smtdv_lib_utils.sv"
`include "smtdv_sequence.sv"
`include "smtdv_sequence_item.sv"
`include "smtdv_component.sv"
`include "smtdv_cfg.sv"
`include "smtdv_event.sv"
`include "smtdv_thread_handler.sv"
`include "smtdv_sequencer.sv"
`include "smtdv_push_sequencer.sv"
`include "smtdv_driver.sv"
`include "smtdv_push_driver.sv"
`include "smtdv_monitor.sv"
`include "smtdv_agent.sv"
`include "smtdv_scoreboard.sv"
`include "smtdv_env.sv"
`include "smtdv_test.sv"
`include "smtdv_runtime_phases.svh"
`include "smtdv_report_server.sv"

`endif
