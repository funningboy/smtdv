
`ifndef __APB_SLAVE_SEQS_CB_SV__
`define __APB_SLAVE_SEQS_CB_SV__




`endif // end of __APB_SLAVE_SEQS_CB_SV__

