`ifndef __SMTDV_TEST_LIST_SV__
`define __SMTDV_TEST_LIST_SV__

  import smtdv_sqlite3_pkg::*;
  import smtdv_stl_pkg::*;

`include "smtdv_base_unittest.sv"

`endif // end of __SMTDV_TEST_LIST_SV__
