
`ifndef __APB_TEST_LIST_SV__
`define __APB_TEST_LIST_SV__

`timescale 1ns/10ps

package test_apb_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import smtdv_sqlite3_pkg::*;
  import smtdv_stl_pkg::*;

  import smtdv_common_pkg::*;
  `include "smtdv_macros.svh"

  `include "apb_defines.svh"
  import apb_pkg::*;
  import apb_seq_pkg::*;

`include "apb_base_test.sv"
`include "apb_setup_test.sv"
`include "apb_rand_test.sv"
`include "apb_stl_test.sv"
`include "apb_retry_test.sv"
`include "apb_err_inject_test.sv"
`include "apb_hijack_test.sv"
`include "apb_polling_test.sv"
`include "apb_interrupt_test.sv"
//`include "apb_fw_ctl_test.sv"
`include "apb_csim_test.sv"

endpackage

`endif // end of __APB_TEST_LIST_SV__
