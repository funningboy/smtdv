../../../../../../../adapters/uvm_sv/uvm_ml_adapter.sv