
`ifndef __XBUS_SLAVE_SEQS_LIB_SV__
`define __XBUS_SLAVE_SEQS_LIB_SV__

`include "xbus_slave_seqs.sv"

`endif
