

virtual class smtdv_scoreboard_cb
  extends
    uvm_callback;
