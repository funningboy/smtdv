uvm_ml_adapter.sv