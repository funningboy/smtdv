uvm_ml_adapter_imp.sv