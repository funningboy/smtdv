
`ifndef __XBUS_SLAVE_SEQS_CB_SV__
`define __XBUS_SLAVE_SEQS_CB_SV__




`endif // end of __XBUS_SLAVE_SEQS_CB_SV__

