// ringbuffer circlebuffer
