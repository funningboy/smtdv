
`ifndef __SMTDV_SLAVE_VSEQS_LIB_SV__
`define __SMTDV_SLAVE_VSEQS_LIB_SV__

`include "smtdv_slave_base_vseq.sv"

`endif // __SMTDV_SLAVE_VSEQS_LIB_SV__
