
//class smtdv_top_graph_builder
//  ) extends
//    smtdv_component#(uvm_env);
//
//  typedef struct
//
//
//endclass : smtdv_top_graph_builder
