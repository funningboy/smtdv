// apb 2 ahb adaptor
