
`ifndef __APB_MASTER_SEQS_LIB_SV__
`define __APB_MASTER_SEQS_LIB_SV__

`include "apb_master_base_seq.sv"
`include "apb_master_atomic_seqs.sv"
`include "apb_master_stl_seq.sv"
`include "apb_master_cfg_seq.sv"
`include "apb_master_irq_seq.sv"

`endif // end of __APB_MASTER_SEQS_LIB_SV__
