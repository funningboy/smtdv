
`ifndef __SMTDV_SQLITE3_PKG_SV__
`define __SMTDV_SQLITE3_PKG_SV__

package smtdv_sqlite3_pkg;
  `include "dpi_smtdv_sqlite3.sv"
endpackage
`endif
