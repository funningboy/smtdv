// cosim with c/systemc
