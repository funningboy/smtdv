
`ifndef __SMTDV_LIB_ALGORITHM_SV__
`define __SMTDV_LIB_ALGORITHM_SV__

`include "smtdv_base_algorithm.sv"
//`inclide "stmtdv_dfs_alg.sv"
//`include "smtdv_scc_alg.sv"

`endif // __SMTDV_LIB_ALGORITHM_SV__
