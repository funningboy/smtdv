// virtual arbiter ...

