../../../../../../../adapters/uvm_sv/uvm_ml_phase.svh