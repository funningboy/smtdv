../../../../../../../adapters/uvm_sv/uvm_ml_tlm1.svh