
// adaptor: extract from sqlite3 db or TLM1 systemc analysis port
`ifndef __XBUS_MASTER_SEQS_CB_SV__
`define __XBUS_MASTER_SEQS_CB_SV__


`endif // __XBUS_MASTER_SEQS_CB_SV__
