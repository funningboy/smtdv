//lock sequence while some block sequence has been asserted
