
`ifndef __CDN_BUSMATRIX_ENV_SV__
`define __CDN_BUSMATRIX_ENV_SV__


`endif // __CDN_BUSMATRIX_ENV_SV__
