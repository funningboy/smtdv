../../../../../../../adapters/uvm_sv/uvm_ml_common.svh