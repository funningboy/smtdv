`ifndef __CDN_BUSMATRIX_SLAVE_VSEQS_LIB_SV__
`define __CDN_BUSMATRIX_SLAVE_VSEQS_LIB_SV__

`include "cdn_slave_base_vseq.sv"

`endif //__CDN_BUSMATRIX_SLAVE_VSEQS_LIB_SV__

