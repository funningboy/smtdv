`ifndef __UART_TEST_LIST_SV__
`define __UART_TEST_LIST_SV__

  import smtdv_sqlite3_pkg::*;

`include "uart_base_test.sv"
`include "uart_seq_test.sv"
//`include "uart_1w1r_test.sv"
//`include "uart_rand_test.sv"
//`include "uart_stl_test.sv"
//`include "uart_err_handle_test.sv"

`endif // end of __UART_TEST_LIST_SV__
