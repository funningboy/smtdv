
`ifndef __DPI_XBUS_IMPORT_SV__
`define __DPI_XBUS_IMPORT_SV__

  import "DPI-C" function chandle dpi_xbus_create_event();

`endif // end of __DPI_XBUS_IMPORT_SV__
