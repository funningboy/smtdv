../../../../../../../adapters/uvm_sv/uvm_ml_hierarchy.svh