`ifndef __APB_MASTER_FW_CTL_VSEQ_SV__
`define __APB_MASTER_FW_CTL_VSEQ_SV__

//class


`endif // __APB_MASTER_FW_CTL_VSEQ_SV__
