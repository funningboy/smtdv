`ifndef __AHB_TEST_LIST_SV__
`define __AHB_TEST_LIST_SV__

`include "ahb_base_env.sv"
`include "ahb_base_test.sv"
`include "ahb_setup_test.sv"
`include "ahb_rand_test.sv"
`include "ahb_stl_test.sv"
`include "ahb_busy_test.sv"
`include "ahb_split_test.sv"
`include "ahb_retry_test.sv"
`include "ahb_err_inject_test.sv"
`include "ahb_hijack_test.sv"
`include "ahb_polling_test.sv"
`include "ahb_interrupt_test.sv"
`include "ahb_incr_test.sv"
`include "ahb_swap_test.sv"
`include "ahb_wrap_test.sv"
`include "ahb_cfg_label_test.sv"
//`include "ahb_fw_ctl_test.sv"
//`include "ahb_csim_test.sv"

`endif // __AHB_TEST_LIST_SV__
