
// cb to TLM2 socket virtual interface
//class
