`ifndef __APB_PKG_SV__
`define __APB_PKG_SV__

package apb_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import smtdv_common_pkg::*;
  `include "smtdv_macros.svh"

  import smtdv_sqlite3_pkg::*;

  import smtdv_stl_pkg::*;

  `include "apb_typedefs.svh"
  `include "apb_item.sv"

  `include "apb_monitor_threads.sv"
  `include "apb_monitor.sv"

  `include "apb_master_cfg.sv"
  `include "apb_master_driver_threads.sv"
  `include "apb_master_driver.sv"
  `include "apb_master_sequencer.sv"
  `include "../seq/apb_master_seqs_lib.sv"
  `include "apb_master_agent.sv"

  `include "apb_slave_cfg.sv"
  `include "apb_slave_driver_threads.sv"
  `include "apb_slave_driver.sv"
  `include "apb_slave_sequencer.sv"
  `include "../seq/apb_slave_seqs_lib.sv"
  `include "apb_slave_agent.sv"

  `include "apb_backdoor.sv"
  `include "apb_scoreboard_threads.sv"
  `include "apb_scoreboard.sv"
  `include "apb_env.sv"
  `include "apb_reg_adapter.sv"
endpackage

`include "apb_if.sv"

`endif
