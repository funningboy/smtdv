`ifndef __AHB_MASTER_SEQS_LIB_SV__
`define __AHB_MASTER_SEQS_LIB_SV__

`include "ahb_master_seqs.sv"
`include "ahb_master_seqs_cb.sv"

`endif // end of __AHB_MASTER_SEQS_LIB_SV__
