
`ifndef __AHB_SLAVE_SEQS_LIB_SV__
`define __AHB_SLAVE_SEQS_LIB_SV__

`include "ahb_slave_base_seq.sv"
`include "ahb_slave_atomic_seqs.sv"
`include "ahb_slave_err_inject_seq.sv"
`include "ahb_slave_hijack_seq.sv"

`endif // __AHB_SLAVE_SEQS_LIB_SV__
