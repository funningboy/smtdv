
`ifndef __SMTDV_UTIL_PKG_SV__
`define __SMTDV_UTIL_PKG_SV__

package smtdv_util_pkg;
  `include "dpi_smtdv_util.sv"
endpackage

`endif // __SMTDV_UTIL_PKG_SV__
