// system look up table as eq idesign spec definition
// [] hash table init
