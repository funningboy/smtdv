`ifndef __AHB_TEST_PKG_SV__
`define __AHB_TEST_PKG_SV__

`timescale 1ns/10ps

package test_ahb_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import smtdv_sqlite3_pkg::*;
  import smtdv_stl_pkg::*;

  import smtdv_common_pkg::*;
  `include "smtdv_macros.svh"

  `include "ahb_defines.svh"
  `include "ahb_macros.svh"

  import ahb_pkg::*;
  import ahb_seq_pkg::*;
  import ahb_vseq_pkg::*;

  `include "ahb_test_lib.sv"

endpackage : test_ahb_pkg

`endif // end of __AHB_TEST_PKG_SV__
