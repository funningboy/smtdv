
`ifndef __CDN_BUSMATRIX_TEST_LIST_SV__
`define __CDN_BUSMATRIX_TEST_LIST_SV__

`include "cdn_busmatrix_env.sv"
`include "cdn_busmatrix_base_test.sv"
`include "cdn_busmatrix_setup_test.sv"

`endif // __CDN_BUSMATRIX_TEST_LIST_SV__

