
`ifndef __SMTDV_LIB_GRAPH_SV__
`define __SMTDV_LIB_GRAPH_SV__

`include "smtdv_attr.sv"
`include "smtdv_node.sv"
`include "smtdv_cmp_node.sv"
`include "smtdv_seq_node.sv"
`include "smtdv_edge.sv"
`include "smtdv_cmp_edge.sv"
`include "smtdv_seq_edge.sv"
`include "smtdv_graph.sv"
`include "smtdv_cmp_graph.sv"
`include "smtdv_seq_graph.sv"

`include "smtdv_seq_graph_builder.sv"
//`include "smtdv_seq_graph_scheduler.sv"
`include "smtdv_cmp_graph_builder.sv"
`include "smtdv_cmp_graph_scheduler.sv"
`include "smtdv_cmp_env.sv"
`include "smtdv_seq_env.sv"

`include "algorithm/smtdv_lib_algorithm.sv"

`endif // __SMTDV_LIB_GRAPH_SV__

