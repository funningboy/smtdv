// about license
