// group model
// register(group)
// order(), sort(),
