
`ifndef __AHB_SLAVE_SEQS_LIB_SV__
`define __AHB_SLAVE_SEQS_LIB_SV__

`include "ahb_slave_seqs.sv"
`include "ahb_slave_seqs_cb.sv"

`endif
