//lock sequence while some block sequence has been asserted

`ifndef __APB_MASTER_MUTEX_VSEQ_SV__
`define __APB_MASTER_MUTRX_VSEQ_SV__

//class apb_master_mutex_vseq
//
//endclass : apb_master_mutex_vseq

`endif // __APB_MASTER_MUTRX_VSEQ_SV__
