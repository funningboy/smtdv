`ifndef __UART_CTRL_TEST_LIST_SV__
`define __UART_CTRL_TEST_LIST_SV__

`endif // end of __UART_CTRL_TEST_LIST_SV__
