// cosim test systemc/c/uvm/v ....
