
//`ifndef __CDN_CPU

