
`ifndef __CDN_TYPEDEFS_SV__
`define __CDN_TYPEDEFS_SV__

`include "bm_params.v"

`endif // __CDN_TYPEDEFS_SV__
