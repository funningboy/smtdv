
`ifndef __AHB_SLAVE_VSEQS_LIB_SV__
`define __AHB_SLAVE_VSEQS_LIB_SV__

`include "ahb_slave_base_vseq.sv"

`endif //__AHB_SLAVE_VSEQS_LIB_SV__

