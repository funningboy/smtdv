`ifndef __AHB_LOCK_WRAP_TEST_SV__
`define __AHB_LOCK_WRAP_TEST_SV__



`endif // end of __AHB_LOCK_WRAP_TEST_SV__
