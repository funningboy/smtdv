//----------------------------------------------------------------------
//   Copyright 2012 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

`ifndef UVM_ML_MACROS_SVH
`define UVM_ML_MACROS_SVH

`define UVM_ML_CONFIG_DB_IMP(T) \
 uvm_config_db_implementation_t #(T)::type_id::set_type_override(uvm_ml_adapter_imp::uvm_ml_singular_config_db_implementation_t #(T)::get_type()); \
 uvm_config_db_implementation_t #(T)::set_imp();

`endif // UVM_ML_MACROS_SVH