// group model
