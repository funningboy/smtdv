`define UVM_KIT_VERSION 13.20-p001
`define UVM_KIT_DATE 2014-01-08
