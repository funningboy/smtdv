// virtual decoder
