
`ifndef __AHB_SLAVE_ATOMIC_SEQS_SV__
`define __AHB_SLAVE_ATOMIC_SEQS_SV__


`endif // end of __AHB_SLAVE_ATOMIC_SEQS_SV__
