// define global/local lookup table to turn on/off each smtdv module
// ex:
//  | path | CPU |  DMA | DDR
// ===========================
//    0    |  0 |    1  | 2
//    1    |  x |    0  | 1
