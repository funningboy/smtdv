

`ifndef __SMTDV_FORCE_VIF_LABEL_SV__
`define __SMTDV_FORCE_VIF_LABEL_SV__

`endif // __SMTDV_FORCE_VIF_LABEL_SV__

