../../../../../../../adapters/uvm_sv/uvm_ml_event.svh