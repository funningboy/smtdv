
`ifndef __SMTDV_SLAVE_SEQS_LIB_SV__
`define __SMTDV_SLAVE_SEQS_LIB_SV__

`include "smtdv_slave_base_seq.sv"
`include "smtdv_slave_fifo_seq.sv"
`include "smtdv_slave_mem_seq.sv"
`include "smtdv_slave_test_seq.sv"

`endif // __SMTDV_SLAVE_SEQS_LIB_SV__
