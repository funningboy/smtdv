
`ifndef __CDN_VIRTUAL_SEQUENCER__
`define __CDN_VIRTUAL_SEQUENCER__
`endif //

