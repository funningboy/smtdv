
// adaptor: extract from sqlite3 db or TLM1 systemc analysis port

`ifndef __XBUS_SLAVE_SEQS_CB_SV__
`define __XBUS_SLAVE_SEQS_CB_SV__

`endif // end of __XBUS_SLAVE_SEQS_CB_SV__

