
`ifndef __AHB_INCR_TEST_SV__
`define __AHB_INCR_TEST_SV__

class ahb_lock_incr_test;

endclass

`endif // end of __AHB_LOCK_INCR_TEST_SV__
