// handle all handler
