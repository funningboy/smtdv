
//`ifndef __SMTDV_EVNET_HANDLER_SV__
//`define __SMTDV_EVENT_HANDLER_SV__
//
//class smtdv_event_handler #
//  extends smtdv_component#(uvm_component);
//
//  bit has_on = 1;
//  longint uuid = -1;
//
//  smtdv_run_event event_q[$];
//
//
//`endif // end of __SMTDV_EVENT_HANDLER_SV__
