
`ifndef __SMTDV_SCOREBOARD_CB_SV__
`define __SMTDV_SCOREBOARD_CB_SV__

/**
* smtdv_scoreboard_cb
*
* @class smtdv_scoreboard_cb
*
*/
class smtdv_scoreboard_cb
  extends
    uvm_object;

endclass : smtdv_scoreboard_cb

`endif // __SMTDV_SCOREBOARD_CB_SV__
