../../../../../../../adapters/uvm_sv/uvm_ml_barrier.svh