
`ifndef __SMTDV_LABEL_HANDLER_SV__
`define __SMTDV_LABEL_HANDLER_SV__

// static handler
class smtdv_label_handler #(
  )extends
  uvm_object;

  bit has_on = 1;
  longint uuid = -1;

  //static
endclass : smtdv_label_handler


`endif // end of __SMTDV_LABEL_HANDLER_SV__
