
`ifndef __APB_SLAVE_SEQS_LIB_SV__
`define __APB_SLAVE_SEQS_LIB_SV__

`include "apb_slave_seqs.sv"
`include "apb_slave_seqs_cb.sv"

`endif
