

`ifndef __SMTDV_UTIL__
`define __SMTDV_UTIL__

  import "DPI-C" function void dpi_getenv(string ienv);
  import "DPI-C" function void dpi_senenv(string ienv, ival);

`endif // __SMTDV_UTIL__
