
`ifndef __CDN_BUSMATRIX_TEST_LIST_SV__
`define __CDN_BUSMATRIX_TEST_LIST_SV__

`include "cdn_base_test.sv"
`include "cdn_setup_test.sv"

`endif // __CDN_BUSMATRIX_TEST_LIST_SV__

