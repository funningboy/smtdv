
`ifndef __UART_CRTL_PKG_SV__
`define __UART_CRTL_PKG_SV__

package uart_ctrl_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import smtdv_common_pkg::*;
  `include "smtdv_macros.svh"

  import smtdv_sqlite3_pkg::*;
  import smtdv_stl_pkg::*;

  import apb_pkg::*;
  import uart_pkg::*;

  `include "uart_ctrl_typedefs.svh"

  `include "uart_ctrl_config.sv"
  `include "uart_ctrl_reg_model.sv"
  `include "uart_apb_s.sv"
  `include "uart_uart_rx.sv"
  `include "uart_uart_tx.sv"
  `include "uart_ctrl_scoreboard.sv"
  `include "uart_ctrl_monitor.sv"
  `include "uart_ctrl_reg_sequencer.sv"
  `include "uart_ctrl_virtual_sequencer.sv"
  `include "uart_ctrl_env.sv"

endpackage : uart_ctrl_pkg

`endif //end of __UART_CTRL_PKG_SV__
