
`ifndef __APB_MASTER_VSEQS_LIB_SV__
`define __APB_MASTER_VSEQS_LIB_SV__

`include "apb_master_base_vseq.sv"
`include "apb_master_1w1r_vseq.sv"
`include "apb_master_stl_vseq.sv"
`include "apb_master_interrupt_vseq.sv"
`include "apb_master_rand_vseq.sv"
`include "apb_master_reset_vseq.sv"

`include "apb_master_retry_vseq.sv"
`include "apb_master_polling_vseq.sv"
`include "apb_master_mutex_vseq.sv"
`include "apb_master_fw_ctl_vseq.sv"
//`include "apb_master_reg_cfg_vseq.sv"

`endif // __APB_MASTER_VSEQS_LIB_SV__
