../../../../../../../adapters/uvm_sv/uvm_ml_phase_service.svh