../../../../../../../adapters/uvm_sv/uvm_ml_serial.svh