
`ifndef __SMTDV_SCOREBOARD_CB_SV__
`define __SMTDV_SCOREBOARD_CB_SV__

class smtdv_scoreboard_cb
  extends
    uvm_object;

endclass

`endif // __SMTDV_SCOREBOARD_CB_SV__
