../../../../../../../adapters/uvm_sv/uvm_ml_resource.svh