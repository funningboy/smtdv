`ifndef __CDN_BUSMATRIX_VSEQS_LIB_SV__
`define __CDN_BUSMATRIX_VSEQS_LIB_SV__

`include "cdn_master_stl_vseq.sv"

`endif // __CDN_BUSMATRIX_VSEQS_LIB_SV__
