
`ifndef __XBUS_TEST_LIST_SV__
`define __XBUS_TEST_LIST_SV__

  import smtdv_sqlite3_pkg::*;
  `include "smtdv_sqlite3_pkg.sv"

`include "xbus_base_test.sv"
`include "xbus_1w1r_test.sv"
`include "xbus_rand_test.sv"

`endif // end of __XBUS_TEST_LIST_SV__
