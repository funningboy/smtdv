../../../../../../../adapters/uvm_sv/uvm_ml_export_dpi.svh