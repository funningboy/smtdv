// about license
// author,
// mail
//
