`ifndef __UART_TX_SEQS_LIB_SV__
`define __UART_TX_SEQS_LIB_SV__

`include "uart_base_seqs.sv"
`include "uart_tx_seqs.sv"
`include "uart_tx_seqs_ref.sv"
`include "uart_tx_seqs_cb.sv"

`endif // __UART_TX_SEQS_LIB_SV__
