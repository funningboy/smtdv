
// adaptor: extract from sqlite3 db or TLM1 systemc analysis channel

