`ifndef __SMTDV_SYSTEM_TABLE_SVH__
`define __SMTDV_SYSTEM_TABLE_SVH__

`endif // __SMTDV_SYSTEM_TABLE_SVH__
