../../../../../../../adapters/uvm_sv/uvm_ml_import_dpi.svh