../../../../../../../adapters/uvm_sv/uvm_ml_blocking_helper.svh