`ifndef __UART_RX_SEQS_LIB_SV__
`define __UART_RX_SEQS_LIB_SV__

`include "uart_rx_base_seq.sv"
`include "uart_rx_seqs_cb.sv"

`endif // __UART_RX_SEQS_LIB_SV__
