
`ifndef __APB_MASTER_SEQS_LIB_SV__
`define __APB_MASTER_SEQS_LIB_SV__

`include "apb_master_seqs.sv"
`include "apb_master_seqs_ref.sv"
`include "apb_master_seqs_cb.sv"

`endif // end of __APB_MASTER_SEQS_LIB_SV__
