
`ifndef __SMTDV_STL_PKG_SV__
`define __SMTDV_STL_PKG_SV__

package smtdv_stl_pkg;
  `include "dpi_smtdv_stl.sv"
endpackage
`endif
