../../../../../../../adapters/uvm_sv/uvm_ml_tlm2.svh