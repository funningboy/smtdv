
`ifndef __APB_TEST_LIST_SV__
`define __APB_TEST_LIST_SV__

  import smtdv_sqlite3_pkg::*;

`include "apb_base_test.sv"
`include "apb_1w1r_test.sv"
`include "apb_rand_test.sv"
`include "apb_stl_test.sv"
`include "apb_err_inject_test.sv"
`include "apb_hijack_test.sv"
`include "apb_csim_test.sv"

`endif // end of __APB_TEST_LIST_SV__
