// not yet implement
