
// adaptor: extract from sqlite3 db / or

