`ifndef __AHB_MASTER_SEQS_LIB_SV__
`define __AHB_MASTER_SEQS_LIB_SV__

`include "ahb_master_base_seq.sv"
`include "ahb_master_atomic_seqs.sv"
`include "ahb_master_stl_seq.sv"
`include "ahb_master_cfg_seq.sv"

`endif // end of __AHB_MASTER_SEQS_LIB_SV__
