
`ifndef __AHB_INTERRUPT_TEST_SV__
`define __AHB_INTERRUPT_TEST_SV__

class apb_interrupt_test
  extends
  apb_base_test;



endclass : apb_interrupt_test

`endif // __AHB_INTERRUPT_TEST_SV__

