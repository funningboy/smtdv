
`ifndef __SMTDV_MASTER_VSEQS_LIB_SV__
`define __SMTDV_MASTER_VSEQS_LIB_SV__

`include "smtdv_master_base_vseq.sv"
`include "smtdv_master_test_vseq.sv"

`endif // __SMTDV_MASTER_VSEQS_LIB_SV__
