
`ifndef __XBUS_MASTER_SEQS_LIB_SV__
`define __XBUS_MASTER_SEQS_LIB_SV__

`include "xbus_master_seqs.sv"
`include "xbus_master_seqs_cb.sv"

`endif // end of __XBUS_MASTER_SEQS_LIB_SV__
