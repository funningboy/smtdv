
`ifndef __SMTDV_SEQ_EDGE_SV__
`define __SMTDV_SEQ_EDGE_SV__

//TODO
`endif // __SMTDV_SEQ_EDGE_SV__
