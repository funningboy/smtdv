
`ifndef __AHB_TEST_LIST_SV__
`define __AHB_TEST_LIST_SV__

  import smtdv_sqlite3_pkg::*;

`include "ahb_base_test.sv"
`include "ahb_lock_incr_test.sv"
`include "ahb_lock_wrap_test.sv"
`include "ahb_lock_swap_test.sv"
`include "ahb_unlock_incr_test.sv"
`include "ahb_unlock_wrap_test.sv"

//`include "ahb_err_handle_test.sv"

`endif // end of __AHB_TEST_LIST_SV__
