
`ifndef __CDN_SRAM_S1_SV__
`define __CDN_SRAM_S1_SV__

class cdn_sram_s1_cfg
  extends
  ahb_slave_cfg

  typedef cdn_sram_s1_cfg cfg_t;

  `uvm_object_param_utils_begin(cfg_t)
  `uvm_object_utils_end

  function new(string name = "cdn_sram_s1_cfg",  smtdv_component cmp=null);
    super.new(name, cmp);
  endfunction : new

endclass : cdn_sram_s1_cfg


class cdn_sram_s1_agent#(
  ADDR_WIDTH = 14,
  DATA_WIDTH = 32)
  extends
  ahb_slave_agent#(
    .ADDR_WIDTH(ADDR_WIDTH),
    .DATA_WIDTH(DATA_WIDTH)
  );

  typedef cdn_sram_s1_agent#(ADDR_WIDTH, DATA_WIDTH) agent_t;

  `uvm_component_param_utils_begin(agent_t)
  `uvm_component_utils_end

  function new(string name = "cdn_sram_s1_agent", uvm_component parent=null);
    super.new(name, parent);
  endfunction : new

endclass : cdn_sram_s1_agent


`endif // __CDN_SRAM_S1_SV__
