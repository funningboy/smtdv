
`ifndef __SMTDV_CIRCULAR_GRAPH_TEST_SV__
`define __SMTDV_CIRCULAR_GRAPH_TEST_SV__

// typedef class smtdv_graph
// typedef class smtdv_node;
// typedef class smtdv_edge;

`endif //__SMTDV_CIRCULAR_GRAPH_TEST_SV__
