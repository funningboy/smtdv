
`ifndef __AHB_INCR_TEST_SV__
`define __AHB_INCR_TEST_SV__

`endif // end of __AHB_LOCK_INCR_TEST_SV__
