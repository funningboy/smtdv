
// convert uart item to other protocol items
