
`ifndef __AHB_SEQ_PKG_SV__
`define __AHB_SEQ_PKG_SV__

`timescale 1ns/10ps

package ahb_seq_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import smtdv_stl_pkg::*;
  import smtdv_sqlite3_pkg::*;

  import smtdv_common_pkg::*;
  import smtdv_common_seq_pkg::*;
  `include "smtdv_macros.svh"

 `include "ahb_defines.svh"
  import ahb_pkg::*;

  `include "ahb_master_seqs_lib.sv"
  `include "ahb_slave_seqs_lib.sv"

endpackage : ahb_seq_pkg

`endif // __AHB_SEQ_PKG_SV__
