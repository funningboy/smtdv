`ifndef __UART_UART_RX_SV__
`define __UART_UART_RX_SV__

